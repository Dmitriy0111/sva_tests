`define ASSERTS_SV