/*
*  File            :   ahb_driver.sv
*  Autor           :   Vlasov D.V.
*  Data            :   2019.11.01
*  Language        :   SystemVerilog
*  Description     :   This is ahb driver
*  Copyright(c)    :   2019 Vlasov D.V.
*/

package test_pkg;

    `include    "classes/ahb_trans.sv"
    `include    "classes/socket.sv"
    `include    "classes/ahb_driver.sv"
    `include    "classes/ahb_monitor.sv"
    `include    "classes/ahb_coverage.sv"
    `include    "classes/base_gen.sv"
    `include    "classes/random_gen.sv"
    `include    "classes/direct_gen.sv"

    `include    "classes/base_test.sv"
    `include    "classes/rand_test.sv"
    `include    "classes/direct_test.sv"
    
endpackage : test_pkg
